asm/test_rom_2.vhd